module Wire( input in, output out );
    assign out=in;
endmodule
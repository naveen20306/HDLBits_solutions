module notgate( input in, output out ); // Declares a module for a NOT gate.
assign out = ~in; // Assigns the inverted value of 'in' to 'out'.
endmodule // Ends the module definition.